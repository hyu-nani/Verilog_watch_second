/* module	date	(
						clk,
						rst,
						);
						
						

	always @ (posedg */